`define COUNT 5
